
class dio_config extends uvm_object;

    `uvm_object_utils(dio_config)

    function new (string name = "");
        super.new(name);
    endfunction : new

endclass : dio_config