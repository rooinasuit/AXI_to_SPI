package clock_pkg;

    `include "clock_driver.sv"
    `include "clock_seq_item.sv"
    `include "clock_sequencer.sv"
    `include "clock_sequences.sv"

endpackage : clock_pkg