package top_pkg;

    `include "test.sv"

endpackage : top_pkg