package test_pkg;

    `include "environment.sv"
    `include "test_base_sequence.sv"
    `include "test_seq_lib.sv"

endpackage : test_pkg