package agents_pkg;

    `include "clock_agent.sv"
    `include "dio_agent.sv"
    `include "spi_slave_agent.sv"

endpackage : agents_pkg