package dio_pkg;

    `include "dio_seq_item.sv"
    `include "dio_sequences.sv"
    `include "dio_sequencer.sv"
    `include "dio_driver.sv"
    `include "dio_monitor.sv"

endpackage : dio_pkg