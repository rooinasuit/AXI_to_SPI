package env_pkg;

`include "virtual_sequencer.sv"
`include "test_sequences.sv"

endpackage : env_pkg