package test_pkg;

    `include "environment.sv"
    `include "test_sequences.sv"

endpackage : test_pkg