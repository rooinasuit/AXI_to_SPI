package macro_pkg;

    `include "monitor_macros.sv"

endpackage : macro_pkg