
class test_sequence_1 extends test_base_sequence;

    `uvm_object_utils(test_sequence_1)

endclass : test_sequence_1 