package dio_seq_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    //
    import dio_pkg::*;
    //
    `include "dio_base_sequence.sv"
    `include "dio_drive_sequence.sv"
    // `include "dio_drive_random_sequence.sv"

endpackage : dio_seq_pkg