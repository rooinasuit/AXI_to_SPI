
class scoreboard_config extends uvm_object;

    `uvm_object_utils(scoreboard_config)

    function new (string name = "scoreaboard_config");
        super.new(name);
    endfunction : new

endclass : scoreboard_config