
interface clock_interface();

    // GLOBAL INPUT SIGNALS
    bit GCLK;

endinterface : clock_interface