package scb_pkg;

    `include "checker.sv"
    `include "ref_model.sv"
    `include "scoreboard.sv"

endpackage : scb_pkg