package clock_seq_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    //
    import clock_pkg::*;
    //
    `include "clock_base_sequence.sv"
    `include "clock_period_sequence.sv"
    `include "clock_state_sequence.sv"

endpackage : clock_seq_pkg