package dio_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    //
    `include "dio_defines.sv"
    //
    `include "dio_config.sv"
    //
    `include "dio_seq_item.sv"
    //
    `include "dio_sequencer.sv"
    `include "dio_driver.sv"
    `include "dio_monitor.sv"
    `include "dio_agent.sv"

endpackage : dio_pkg