package test_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import env_pkg::*;

    `include "test_base_sequence.sv"
    `include "test_seq_lib.sv"
    `include "test.sv"

endpackage : test_pkg