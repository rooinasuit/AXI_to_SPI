package seq_pkg;

`include "virtual_sequencer.sv"
`include "test_sequences.sv"

endpackage : seq_pkg