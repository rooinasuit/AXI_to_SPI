`define CHECKER_DECLARE() \

`define CHECKER_CREATE() \
