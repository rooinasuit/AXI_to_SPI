
interface clk_interface();

    // GLOBAL INPUT SIGNALS
    bit GCLK;

endinterface : clk_interface