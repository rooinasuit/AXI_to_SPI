package top_pkg;

    `include "test_sequences.sv"
    `include "test.sv"

endpackage : top_pkg