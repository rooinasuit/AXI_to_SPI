
class clock_config extends uvm_object;

    `uvm_object_utils(clock_config)

    function new (string name = "");
        super.new(name);
    endfunction : new

endclass : clock_config