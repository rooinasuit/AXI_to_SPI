package scb_pkg;

    `include "checker.sv"
    `include "ref_model.sv"

endpackage : scb_pkg