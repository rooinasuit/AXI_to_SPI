package clock_pkg;

    `include "clock_seq_item.sv"
    `include "clock_base_sequence.sv"
    `include "clock_seq_lib.sv"
    `include "clock_sequencer.sv"
    `include "clock_driver.sv"

endpackage : clock_pkg