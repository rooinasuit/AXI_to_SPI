
interface clock_interface();

    // GLOBAL INPUT SIGNALS
    logic GCLK;

endinterface : clock_interface